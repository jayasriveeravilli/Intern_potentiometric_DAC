* C:\Users\drsur\Documents\LTspiceXVII\10bit.asc
XX3 N001 o10 a9 N004 switch
R1 N002 N003 0.625k
XX1 a0 a1 a2 a3 a4 a5 a6 a7 a8 N001 ir10 N002 9bit
XX2 a0 a1 a2 a3 a4 a5 a6 a7 a8 N004 N003 or10 9bit
V1 a0 0 PWL(0 0 0.99 0 1 5 1.99 5 2 0 2.99 0 3 5 3.99 5 4 0)
V2 a1 0 PWL(0 0 1.99 0 2 5 2.99 5 3 0 4 0)
V3 0 a2 PWL(0 0 0.99 0 1 5 2.99 5 3 0 4 0)
V4 0 a3 PWL(0 5 0.99 5 1 0 1.99 0 2 5 2.99 5 3 0 4 0)
V5 a8 0 PWL(0 0 1.99 0 2 5 3.99 5 4 0)
V6 a7 0 PWL(0 0 0.99 0 1 5 1.99 5 2 0 4 0)
V7 a6 0 PWL(0 5 0.99 5 1 0 2.99 0 3 5 3.99 5 4 0)
V8 a5 0 PWL(0 5 2.99 5 3 0 4 0)
V9 a4 0 PWL(0 0 0.99 0 1 5 1.99 5 2 0 4 0)
V10 a9 0 PWL(0 0 0.99 0 1 5 3.99 5 4 0)

* block symbol definitions
.subckt switch in1 Vout d_in in2
M1 N001 N004 N003 N001 PMOS
M2 in1 N003 Vout N002 PMOS
M3 Vout d_in in2 Vout PMOS
M4 in1 d_in Vout Vout NMOS
M5 Vout N003 in2 N005 NMOS
M6 N003 N004 0 0 NMOS
V1 N001 0 3.3
.model n_mos NMOS (LEVEL=8 VERSION=3.2 TNOM=27 TOX=4.1E-9 XJ=1E-7 NCH=2.3549E17 VTH0=0.3823463 K1=0.5810697
*+            K2=4.774618E-3 K3=0.0431669 K3B=1.1498346 W0=1E-7 NLX=1.910552E-7 DVT0W=0 DVT1W=0 DVT2W=0
*+            DVT0=1.2894824 DVT1=0.3622063 DVT2=0.0713729 U0=280.633249 UA=-1.208537E-9 UB=2.158625E-18
*+            UC=5.342807E-11 VSAT=9.366802E4 A0=1.7593146 AGS=0.3939741 B0=-6.413949E-9 B1=-1E-7 KETA=-5.180424E-4
*+            A1=0 A2=1 RDSW=105.5517558 PRWG=0.5 PRWB=-0.1998871 WR=1 WINT=7.904732E-10 LINT=1.571424E-8 XL=0
*+            XW=-1E-8 DWG=1.297221E-9 DWB=1.479041E-9 VOFF=-0.0955434 NFACTOR=2.4358891 CIT=0 CDSC=2.4E-4 CDSCD=0
*+            CDSCB=0 ETA0=3.104851E-3 ETAB=-2.512384E-5 DSUB=0.0167075 PCLM=0.8073191 PDIBLC1=0.1666161 PDIBLC2=3.112892E-3
*+            PDIBLCB=-0.1 DROUT=0.7875618 PSCBE1=8E10 PSCBE2=9.213635E-10 PVAG=3.85243E-3 DELTA=0.01 RSH=6.7 MOBMOD=1
*+            PRT=0 UTE=-1.5 KT1=-0.11 KT1L=0 KT2=0.022 UA1=4.31E-9 UB1=-7.61E-18 UC1=-5.6E-11 AT=3.3E4 WL=0 WLN=1
*+            WW=0 WWN=1 WWL=0 LL=0 LLN=1 LW=0 LWN=1 LWL=0 CAPMOD=2 XPART=0.5 CGDO=7.08E-10 CGSO=7.08E-10 CGBO=1E-12
*+            CJ=9.68858E-4 PB=0.8 MJ=0.3864502 CJSW=2.512138E-10 PBSW=0.809286 MJSW=0.1060414 CJSWG=3.3E-10 PBSWG=0.809286
*+            MJSWG=0.1060414 CF=0 PVTH0=-1.192722E-3 PRDSW=-5 PK2=6.450505E-5 WKETA=-4.27294E-4 LKETA=-0.0104078
*+            PU0=6.3268729 PUA=2.226552E-11 PUB=0 PVSAT=969.1480157 PETA0=1E-4 PKETA=-1.049509E-3)
.model p_mos PMOS (LEVEL=8 VERSION=3.2 TNOM=27 TOX=4.1E-9 XJ=1E-7 NCH=4.1589E17 VTH0=-0.3938813 K1=0.5479015
*+            K2=0.0360586 K3=0.0993095 K3B=5.7086622 W0=1E-6 NLX=1.313191E-7 DVT0W=0 DVT1W=0 DVT2W=0 DVT0=0.4911363
*+            DVT1=0.2227356 DVT2=0.1 U0=115.6852975 UA=1.505832E-9 UB=1E-21 UC=-1E-10 VSAT=1.329694E5 A0=1.7590478
*+            AGS=0.3641621 B0=3.427126E-7 B1=1.062928E-6 KETA=0.0134667 A1=0.6859506 A2=0.3506788 RDSW=168.5705677
*+            PRWG=0.5 PRWB=-0.4987371 WR=1 WINT=0 LINT=3.028832E-8 XL=0 XW=-1E-8 DWG=-2.349633E-8 DWB=-7.152486E-9
*+            VOFF=-0.0994037 NFACTOR=1.9424315 CIT=0 CDSC=2.4E-4 CDSCD=0 CDSCB=0 ETA0=0.0608072 ETAB=-0.0426148
*+            DSUB=0.7343015 PCLM=3.2579974 PDIBLC1=7.229527E-6 PDIBLC2=0.025389 PDIBLCB=-1E-3 DROUT=0 PSCBE1=1.454878E10
*+            PSCBE2=4.202027E-9 PVAG=15 DELTA=0.01 RSH=7.8 MOBMOD=1 PRT=0 UTE=-1.5 KT1=-0.11 KT1L=0 KT2=0.022 UA1=4.31E-9
*+            UB1=-7.61E-18 UC1=-5.6E-11 AT=3.3E4 WL=0 WLN=1 WW=0 WWN=1 WWL=0 LL=0 LLN=1 LW=0 LWN=1 LWL=0 CAPMOD=2 XPART=0.5
*+            CGDO=6.32E-10 CGSO=6.32E-10 CGBO=1E-12 CJ=1.172138E-3 PB=0.8421173 MJ=0.4109788 CJSW=2.242609E-10 PBSW=0.8            +            MJSW=0.3752089 CJSWG=4.22E-10 PBSWG=0.8 MJSWG=0.3752089 CF=0 PVTH0=1.888482E-3 PRDSW=11.5315407 PK2=1.559399E-3
*+            WKETA=0.0319301 LKETA=2.955547E-3 PU0=-1.1105313 PUA=-4.62102E-11 PUB=1E-21 PVSAT=50 PETA0=1E-4 PKETA=-4.346368E-3)
.ends switch

.subckt 9bit a0 a1 a2 a3 a4 a5 a6 a7 a8 o9 ir9 or9
XX1 N001 ir9 N002 a0 a1 a2 a3 a4 a5 a6 a7 8bit
XX2 N004 N003 or9 a0 a1 a2 a3 a4 a5 a6 a7 8bit
R1 N002 N003 0.625k
XX3 N001 o9 a8 N004 switch
.ends 9bit

.subckt 8bit o8 ir8 or8 a0 a1 a2 a3 a a5 a6 a7
XX1 N001 ir8 N002 a0 a1 a2 a3 a4 a5 a6 7bit
XX2 N003 P001 or8 a0 a1 a2 a3 a4 a5 a6 7bit
XX3 N001 o8 a7 N003 switch
R1 N002 P001 0.625k
.ends 8bit

.subckt 7bit o7 ir7 or7 a0 a1 a2 a3 a4 a5 a6
XX1 N001 ir7 N002 a0 a1 a2 a3 a4 a5 6bit
XX2 N004 N003 or7 a0 a1 a2 a3 a4 a5 6bit
XX3 N001 o7 a6 N004 switch
R1 N002 N003 0.625k
.ends 7bit

.subckt 6bit o6 ir6 or6 a0 a1 a2 a3 a4 a5
XX1 a0 a1 a2 a3 a4 ir6 N002 N001 5bit
XX2 a0 a1 a2 a3 a4 N003 or6 N004 5bit
R1 N002 N003 0.625k
XX3 N001 o6 a5 N004 switch
.ends 6bit

.subckt 5bit a0 a1 a2 a3 a4 ri5 ro5 o5
XX1 ri5 N002 N001 a0 a1 a2 a3 4bit
XX2 N003 ro5 N004 a0 a1 a2 a3 4bit
XX3 N001 o5 a4 N004 switch
R1 N002 N003 0.625k
.ends 5bit

.subckt 4bit rin r0 o4 a0 a1 a2 a3
XX1 a0 a1 a2 N001 rin N002 3bit
XX2 a0 a1 a2 N004 N003 ro 3bit
XX3 N001 o4 a3 N004 switch
R1 N002 N003 0.625k
.ends 4bit

.subckt 3bit a0 a1 a2 o3 inres outres
XX1 a0 a1 N001 inres P001 2bit
XX2 a0 a1 N003 N002 outres 2bit
XX3 N001 o3 a2 N003 switch
R1 P001 N002 0.625k
.ends 3bit

.subckt 2bit a0 a1 o2 inpin outpin
XX1 inpin N001 a0 N002 switch
XX2 N003 N004 a0 N005 switch
XX3 N001 o2 a1 N004 switch
R1 inpin N002 0.625k
R2 N002 N003 0.625k
R3 N003 N005 0.625k
R4 N005 outpin 0.625k
.ends 2bit

.model NMOS NMOS
.model PMOS PMOS
*.lib C:\Users\drsur\Documents\LTspiceXVII\lib\cmp\standard.mos
* 9b
* 9b
.tran 100ms
*.backanno
.end
